library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CU is
    Port ( 
			  op : in  STD_LOGIC_VECTOR (1 downto 0);
           op3 : in  STD_LOGIC_VECTOR (5 downto 0);
           
           ALUOP : out  STD_LOGIC_VECTOR (5 downto 0));
end CU;

architecture Behavorial of CU is

begin
	
	process(op,op3)
	
	begin
		ALUOP <= "000000";
					if(op = "10")then				
						case op3 is
							when "000000" => -- ADD
								
								ALUOP <= "000000";							
							when "000100"=> --sub
								
								ALUOP <= "000100";							
							when "000001" => --and
								
								ALUOP <= "000001";	
							when "000101" => --andn
								
								ALUOP <= "000101";
							when "000010" => -- or
								
								ALUOP <= "000010";
							when "000110" => -- orn
								
								ALUOP <= "000110";
							when "000011" => -- xor	
								
								ALUOP <= "000011";
							when "000111" => -- xnor
								
								ALUOP <= "000111";
								
							when others => -- Implementar demas instrucciones
								
								ALUOP <= "000000";
						end case;
					else
						ALUOP <= "000000";
						
					end if;
	
	end process;
end Behavorial;